--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:16:09 12/09/2013
-- Design Name:   
-- Module Name:   C:/Users/Madkiche/Desktop/modulador/modulador/tb_modo.vhd
-- Project Name:  modulador
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: modo
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_modo IS
END tb_modo;
 
ARCHITECTURE behavior OF tb_modo IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT modo
    PORT(
         sincro_modo : IN  std_logic;
         clk : IN  std_logic;
         reset : IN  std_logic;
         valor_modo : BUFFER  std_logic_vector(1 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal sincro_modo : std_logic := '0';
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';

 	--Outputs
   signal valor_modo : std_logic_vector(1 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: modo PORT MAP (
          sincro_modo => sincro_modo,
          clk => clk,
          reset => reset,
          valor_modo => valor_modo
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		reset <= '1';
		wait for 43 ns;
		reset <= '0';
      wait for clk_period*10;
		sincro_modo <= '1';
		wait for 85 ns;
		sincro_modo <= '0';
      -- insert stimulus here 

      wait;
   end process;

END;
